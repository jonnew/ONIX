----------------------------------------------------------------------------------
--This is the SPI input module that takes a serial command and make it a parallel sequence
----------------------------------------------------------------------------------
library IEEE;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_1164.ALL;

entity SPI_input is
end SPI_input;

architecture Behavioral of SPI_input is

begin


end Behavioral;

