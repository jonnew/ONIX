// NB: colors.mem was generated using colors.py. There are lots of hard-coded
// constants in here that would need to be changed if the number of colors or
// their order is altered

`include "./ws2811/ws2811.v"

module neopix_controller # (
    parameter CLK_RATE_HZ   = 50_000_000
) (
    // Clock and reset
    input   wire            i_clk,
    input   wire            i_reset,

    // Derived from host to breakout slow word
    input   wire            i_acq_running,
    input   wire            i_acq_reset_done,
    input   wire    [3:0]   i_ledlevel,
    input   wire    [1:0]   i_ledmode,
    input   wire    [1:0]   i_porta_status,
    input   wire    [1:0]   i_portb_status,
    input   wire    [1:0]   i_portc_status,
    input   wire    [1:0]   i_portd_status,
    input   wire    [11:0]  i_aio_dir,
    input   wire    [1:0]   i_harp_conf, // TODO
    input   wire    [15:0]  i_gpio_dir,  // TODO

    // Link power
    input   wire    [3:0]   i_link_pow,

    // HARP heartbeat
    input   wire            i_harp_hb,

    // Button press state
    input   wire    [5:0]   i_button,

    // Digital IO
    input   wire    [7:0]   i_din_state,
    input   wire    [7:0]   i_dout_state,

    // Neopixel control signal
    output  wire            o_neopix

    // Debug
    //output  wire    [7:0]   o_quotient_debug
);

// Colors
reg [23:0] off,
           blue,
           orange,
           green,
           red,
           purple,
           brown ,
           pink ,
           white ,
           yellow,
           cyan;

// This is ultra hardcoded for the particular color set generated by colors.py
reg [23:0] colors [0:159]; //  (1 << $clog2(160)) - 1];
reg [7:0] color_addr;
reg [3:0] color_idx, color_idx_last;
reg [23:0] color;

initial $readmemh("colors.mem", colors);
initial off = 0;

// RAM address
always @ (posedge i_clk) begin

    color_idx_last <= color_idx;

    if (i_reset) begin
        color_addr <= 0;
        color_idx <= 0;
    end else if (color_idx == 0) begin
        color_addr <= 144 + {4'b0000, i_ledlevel};
        color_idx <= 9;
    end else begin
        color_addr <= color_addr - 16;
        color_idx <= color_idx - 1;
    end
end

// RAM access
always @ (posedge i_clk) begin
    color <= colors[color_addr];
end

always @ (posedge i_clk) begin

    case (color_idx_last)
        0:
            blue <= color;
        1:
            orange <= color;
        2:
            green <= color;
        3:
            red <= color;
        4:
            purple <= color;
        5:
            brown <= color;
        6:
            pink <= color;
        7:
            white <= color;
        8:
            yellow <= color;
        9:
            cyan <= color;

    endcase
end

// Neopixel color state
reg [23:0] rgb [0:40];

// LED use levels
reg dark = 1'b0;
reg released = 1'b1;
wire led_mode1 = ~dark & (i_ledmode[0] | i_ledmode[1]);
wire led_mode2 = ~dark & i_ledmode[1];
wire led_mode3 = ~dark & (i_ledmode[0] & i_ledmode[1]);

always @ (posedge i_clk) begin

    if (i_button[0] && released) begin
        dark <= dark + 1;
        released <= 1'b0;
    end else if (!i_button[0]) begin
        released <= 1'b1;
    end
end

// LED color logic
always @ (*) begin

    rgb[0] = led_mode1 ? yellow : off;

    rgb[1] = led_mode2 ?
            (i_acq_reset_done ?
            (i_acq_running ?
            (i_harp_hb ?
            red : off) : red) : purple) : off;

    //rgb[1] = (led_mode3 & i_button[5]) ? blue : off;
    rgb[2] = (led_mode3 & i_button[5]) ? blue : off;
    rgb[3] = (led_mode3 & i_button[4]) ? blue : off;
    rgb[4] = (led_mode3 & i_button[3]) ? blue : off;
    rgb[5] = (led_mode3 & i_button[2]) ? blue : off;
    rgb[6] = (led_mode3 & i_button[1]) ? blue : off;

    rgb[7] = off; // TODO: "Host"
    rgb[8] = (led_mode2 & i_harp_hb) ? red : off;

    rgb[9]  = (led_mode3 & i_din_state[0]) ? green : off;
    rgb[10] = (led_mode3 & i_din_state[1]) ? green : off;
    rgb[11] = (led_mode3 & i_din_state[2]) ? green : off;
    rgb[12] = (led_mode3 & i_din_state[3]) ? green : off;
    rgb[13] = (led_mode3 & i_din_state[4]) ? green : off;
    rgb[14] = (led_mode3 & i_din_state[5]) ? green : off;
    rgb[15] = (led_mode3 & i_din_state[6]) ? green : off;
    rgb[16] = (led_mode3 & i_din_state[7]) ? green : off;

    rgb[17] = (led_mode3 & i_dout_state[7]) ? green : off;
    rgb[18] = (led_mode3 & i_dout_state[6]) ? green : off;
    rgb[19] = (led_mode3 & i_dout_state[5]) ? green : off;
    rgb[20] = (led_mode3 & i_dout_state[4]) ? green : off;
    rgb[21] = (led_mode3 & i_dout_state[3]) ? green : off;
    rgb[22] = (led_mode3 & i_dout_state[2]) ? green : off;
    rgb[23] = (led_mode3 & i_dout_state[1]) ? green : off;
    rgb[24] = (led_mode3 & i_dout_state[0]) ? green : off;

    // Port A (HS3 on the board)
    if (!led_mode1 || i_porta_status == 1)
        rgb[25] = off;
    else if (i_porta_status == 3)
        rgb[25] = i_acq_running ? (i_harp_hb ? red : off) : red;
    else if (i_link_pow[3] && i_porta_status == 2)
        rgb[25] = purple;
    else
        rgb[25] = off;

    // Port B (HS2 on the board)
    if (!led_mode1 || i_portb_status == 1)
        rgb[26] = off;
    else if (i_portb_status == 3)
        rgb[26] = i_acq_running ? (i_harp_hb ? red : off) : red;
    else if (i_link_pow[2] && i_portb_status == 2)
        rgb[26] = purple;
    else
        rgb[26] = off;

    // Port C (HS1 on the board)
    if (!led_mode1 || i_portc_status == 1)
        rgb[27] = off;
    else if (i_portc_status == 3)
        rgb[27] = i_acq_running ? (i_harp_hb ? red : off) : red;
    else if (i_link_pow[1] && i_portc_status == 2)
        rgb[27] = purple;
    else
        rgb[27] = off;

    // Port D (HS0 on the board)
    if (!led_mode1 || i_portd_status == 1)
        rgb[28] = off;
    else if (i_portd_status == 3)
        rgb[28] = i_acq_running ? (i_harp_hb ? red : off) : red;
    else if (i_link_pow[0] && i_portd_status == 2)
        rgb[28] = purple;
    else
        rgb[28] = off;

    // Analog IO
    rgb[29] = led_mode3 ? (i_aio_dir[11] ? cyan : brown) : off;
    rgb[30] = led_mode3 ? (i_aio_dir[10] ? cyan : brown) : off;
    rgb[31] = led_mode3 ? (i_aio_dir[9]  ? cyan : brown) : off;
    rgb[32] = led_mode3 ? (i_aio_dir[8]  ? cyan : brown) : off;
    rgb[33] = led_mode3 ? (i_aio_dir[7]  ? cyan : brown) : off;
    rgb[34] = led_mode3 ? (i_aio_dir[6]  ? cyan : brown) : off;
    rgb[35] = led_mode3 ? (i_aio_dir[0]  ? cyan : brown) : off;
    rgb[36] = led_mode3 ? (i_aio_dir[1]  ? cyan : brown) : off;
    rgb[37] = led_mode3 ? (i_aio_dir[2]  ? cyan : brown) : off;
    rgb[38] = led_mode3 ? (i_aio_dir[3]  ? cyan : brown) : off;
    rgb[39] = led_mode3 ? (i_aio_dir[4]  ? cyan : brown) : off;
    rgb[40] = led_mode3 ? (i_aio_dir[5]  ? cyan : brown) : off;

end

// Currently addressed LED
wire [5:0] led_addr;

// Neopixel control
ws2811 # (
    .NUM_LEDS(41),
    .SYSTEM_CLOCK(CLK_RATE_HZ)
) neopix (
    .clk(i_clk),
    .reset(i_reset),
    .address(led_addr),
    .red_in(rgb[led_addr][23:16]),
    .green_in(rgb[led_addr][15:8]),
    .blue_in(rgb[led_addr][7:0]),
    .DO(o_neopix)
);

endmodule
