// Facts about this design:
//
// 1. It is meant, insofar as possible, to be a zero-latency "view" into the
// hardware on the breakout board that is controlled by the host.
//
// 2. The clock governing the whole board is derived from an LVDS line coming
// from the host board. The PLL is locked to this clock for data transmission.
// Data coming to the breakout board is synchronous to the LVDS clock and
// data going out of the breakout board is sychronous to the PLL-generated
// clock.
//
// 3. Have a look at host_to_breakout.v and breakout_to_host.v for
// descriptions of data packet format.
//
// 4. There is no error correction or CRC, currently.

//`include "pll_10_60.v"
`include "pll_10_60_2ns.v"
//`include "pll_16_60_2ns.v"
//`include "pll_16_60.v"
`include "breakout_to_host.v"
`include "host_to_breakout.v"
`include "user_io.v"
`include "harp_sync.v"
`include "neopix_controller.v"

module breakout (
    input   wire            XTAL,    // 16MHz clock
    input   wire            D_IN0,   // Manual SB_IO means I can't use array
    input   wire            D_IN1,
    input   wire            D_IN2,
    input   wire            D_IN3,
    input   wire            D_IN4,
    input   wire            D_IN5,
    input   wire            D_IN6,
    input   wire            D_IN7,
    output  wire    [7:0]   D_OUT,
    input   wire    [1:0]   LVDS_IN,
    output  wire    [2:0]   LVDS_OUT,
    inout   wire            I2C_SCL,
    inout   wire            I2C_SDA,
    output  wire            HARP_CLK_OUT,
    output  wire            LED,   // User/boot LED next to power LED
    output  wire            USBPU, // USB pull-up resistor
    output  wire            NEOPIX

    //// Simulation
    //output   wire            I2C_SCL,
    //output   wire            I2C_SDA,
    //input   wire             PLL_SIM
);

// Internal nets
reg reset;
wire [5:0] buttons;
wire [3:0] link_pow;

// Host to breakout slow word results
wire [7:0] ledlevel;
wire [1:0] ledmode;
wire [1:0] porta_status;
wire [1:0] portb_status;
wire [1:0] portc_status;
wire [1:0] portd_status;
wire [11:0] aio_dir;
wire [1:0] harp_conf;
wire [15:0] gpio_dir;

// D_INs with pullup applied
wire [7:0] d_in_pu;

// Main system clock
// ---------------------------------------------------------------
wire sys_clk;
wire pll_locked ;

pll_10_60_2ns pll_sys(LVDS_IN[0], sys_clk, pll_locked); // 60 MHz sys clk

// Testing
//pll_16_60 pll_sys(XTAL, sys_clk, pll_locked); // 60 MHz sys clk

// Simulation
//assign reset = 0;
//assign sys_clk = PLL_SIM;

// Power on reset
reg [8:0] reset_cnt = 0;
assign reset = ~reset_cnt[8];
always @(posedge sys_clk)
    if (pll_locked)
        reset_cnt <= reset_cnt + reset;

// IO expander
// ---------------------------------------------------------------

user_io # (
    .CLK_RATE_HZ(60_000_000),
    .I2C_CLK_RATE_HZ(400_000)
) uio (
    .i_clk(sys_clk),
    .i_reset(reset),
    .i_porta_status(porta_status),
    .i_portb_status(portb_status),
    .i_portc_status(portc_status),
    .i_portd_status(portd_status),
    .o_button(buttons),
    .o_link_pow(link_pow),
    .io_scl(I2C_SCL),
    .io_sda(I2C_SDA)
    //.o_state(D_OUT[4:0])
);

// Breakout to host
// ---------------------------------------------------------------
breakout_to_host b2h (
    .i_clk(sys_clk),
    .i_port(D_IN),
    .i_button(buttons),
    .i_link_pow(link_pow),
    .o_clk_s(LVDS_OUT[0]),
    .o_d0_s(LVDS_OUT[1]),
    .o_d1_s(LVDS_OUT[2])
);

// Host to breakout
// ---------------------------------------------------------------
host_to_breakout h2b (
    .i_clk(sys_clk), // Synchronous to LVDS_IN[0]
    .i_clk_s(LVDS_IN[0]),
    .i_d0_s(LVDS_IN[1]),
    .o_port(D_OUT),
    .o_ledlevel(ledlevel),
    .o_ledmode(ledmode),
    .o_porta_status(porta_status),
    .o_portb_status(portb_status),
    .o_portc_status(portc_status),
    .o_portd_status(portd_status),
    .o_aio_dir(aio_dir),
    .o_harp_conf(harp_conf),
    .o_gpio_dir(gpio_dir)
    //.o_slow_valid(slow_word_valid),
    //.o_slow_value(slow_word),
    //.o_reset(open), // TODO
);

// HARP
// ---------------------------------------------------------------
harp_sync # (
    .CLK_RATE_HZ(60_000_000)
) sync (
    .clk(sys_clk),
    .reset(reset),
    .run('b1),
    .TX(HARP_CLK_OUT),
    .LED(harp_hb)
);

// Neopixel control
// ---------------------------------------------------------------
neopix_controller # (
    .CLK_RATE_HZ(60_000_000)
) neopix (
    .i_clk(sys_clk),
    .i_reset(reset),
    .i_harp_hb(harp_hb),
    .i_pll_lock(pll_locked),
    .i_link_pow(link_pow),
    .i_button(buttons),
    .i_din_state(d_in_pu),
    .i_dout_state(D_OUT),
    .i_ledlevel(ledlevel),
    .i_ledmode(ledmode),
    .i_porta_status(porta_status),
    .i_portb_status(portb_status),
    .i_portc_status(portc_status),
    .i_portd_status(portd_status),
    .i_aio_dir(aio_dir),
    .i_harp_conf(harp_conf),
    .i_gpio_dir(gpio_dir),
    .o_neopix(NEOPIX)
);

// IO settings
// ---------------------------------------------------------------

// Ony indicate progrmaming mode
assign LED = 0; //pll_locked;

// Drive USB pull-up resistor to '0' to disable USB
assign USBPU = 0;

// Enable pullups on the digital input port
SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din0 (
  .PACKAGE_PIN(D_IN0),
  .D_IN_0(d_in_pu[0])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din1 (
  .PACKAGE_PIN(D_IN1),
  .D_IN_0(d_in_pu[1])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din2 (
  .PACKAGE_PIN(D_IN2),
  .D_IN_0(d_in_pu[2])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din3 (
  .PACKAGE_PIN(D_IN3),
  .D_IN_0(d_in_pu[3])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din4 (
  .PACKAGE_PIN(D_IN4),
  .D_IN_0(d_in_pu[4])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din5 (
  .PACKAGE_PIN(D_IN5),
  .D_IN_0(d_in_pu[5])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din6 (
  .PACKAGE_PIN(D_IN6),
  .D_IN_0(d_in_pu[6])
);

SB_IO #(
  .PIN_TYPE(6'b 0000_01),
  .PULLUP(1'b 1)
) din7 (
  .PACKAGE_PIN(D_IN7),
  .D_IN_0(d_in_pu[7])
);

endmodule
